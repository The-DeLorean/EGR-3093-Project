----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Dorian Quimby
-- 
-- Create Date: 04/16/2024 04:35:17 PM
-- Design Name: 
-- Module Name: navigation_check - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: This module takes in the location of a game object (Pacman or ghost).
-- It will return flags based on whether certain moves are possible.
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;


-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity navigation_check is
    Port ( x_pos : in integer;
           y_pos : in integer;
           down  : in std_logic;
           --input of map?
           collision : out std_logic
           --right : out std_logic;
           --up : out std_logic;
           --down : out std_logic
           );
end navigation_check;

architecture Behavioral of navigation_check is
constant rom_depth : natural := 448; --32
constant rom_width : natural := 392;--28
signal collision_i : std_logic:='0';

signal wall_bit: std_logic:='0';
signal y_pos_i : integer;
signal x_pos_i : integer;

type wall_type is array (0 to rom_depth -1) of std_logic_vector(rom_width - 1 downto 0);
--origin (124, 5)
constant walls : wall_type :=(
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111100000000000000000000000000001111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000001111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000011111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000011111111111111111111111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

--constant walls : wall_type :=(
--                            "0000000000001100000000000011",
--                            "0111101111101101111101111011",
--                            "0111101111101101111101111011",
--                            "0111101111101101111101111011",
--                            "0000000000000000000000000011",
--                            "0111101101111111101101111011",
--                            "0111101101111111101101111011",
--                            "0000001100001100001100000011",
--                            "1111101111101101111101111111",
--                            "0000101111101101111101000011",
--                            "0000101100000000001101000011",
--                            "0000101101110011101101000011",
--                            "1111101101000000101101111111",
--                            "0000000001000000100000000011",
--                            "1111101101000000101101111111",
--                            "0000101101111111101101000011",
--                            "0000101100000000001101000011",
--                            "0000101101111111101101000011",
--                            "1111101101111111101101111111",
--                            "0000000000001100000000000011",
--                            "0111101111101101111101111011",
--                            "0111101111101101111101111011",
--                            "0001100000000000000001100011",
--                            "1101101101111111101101101111",
--                            "1101101101111111101101101111",
--                            "0000001100001100001100000011",
--                            "0111111111101101111111111011",
--                            "0111111111101101111111111011",
--                            "0000000000000000000000000011",
--                            "1111111111111111111111111111",
--                            "1111111111111111111111111111",
--                            "1111111111111111111111111111");

begin 

process
begin
    if down ='0' then
        wall_bit<=walls(y_pos+13)(x_pos);
        if wall_bit='1' then
            collision_i<='1';
        else 
             collision_i<='0';
        end if;
    end if;
--    if down ='0' then
--        y_pos_i<=y_pos + 1;
--        x_pos_i<=x_pos;
--    end if;
----    for i in 0 to rom_depth - 1 loop 
----        for j in 0 to rom_width - 1 loop
----            wait for 1 ns;
----            --assign wall bit
----            wall_bit <= walls()(j);
            
--           -- if( wall_bit = '1' ) then --if there is actually a block there
----                if( ( abs( (j*14 + 124) - x_pos ) < 50 )
----                AND ( abs( (i*14 + 5) - y_pos ) < 50 ) ) then --if object is nearby
----                    if (    ((y_pos +12 >= (i*14) + 5) And (x_pos >= (j*14)+124 -12 and x_pos<= (j*14)+124+12)) AND down='0' ) then --OR
----                          --  if((y_pos+7<= (i*14) + 5 - 6) OR
------                            (y_pos >= (i*14) + 5 + 6) OR
------                            (x_pos >= (j*14) + 124 + 6) OR
------                            (x_pos+7 <= (j*14) + 124 - 6) ) then --check for collision
----                        collision_i <= '1'; --collision
----                    end if;
----               end if;
----                        --I
----                        if not(x_pos = (j*14)+124 and x_pos+14 = (j*14)+124+14) then
----                            collision_i <= '0'; -- no collision
----                        end if;


----            WORKS BEST I THINK Unccoment lines below to have it almost work perfectly
--    for i in 0 to rom_depth - 1 loop 
--        for j in 0 to rom_width - 1 loop
--            wait for 1 ns;
--            --assign wall bit
--            wall_bit <= walls(i)(j);
--           if( wall_bit = '1' ) then --if there is actually a block there
--                if(down='0') then
--                        if (    ((y_pos_i  >= (i*14) + 6-14) and y_pos_i<(i*14) And x_pos_i >= (j*14)+124 and x_pos_i <= (j*14)+124+14)) then
--                            collision_i<='1'; -- collision
   
--                       end if;
--                end if;
--           end if;
--        end loop;
--    end loop;  
end process;

collision <= collision_i;
end Behavioral;
